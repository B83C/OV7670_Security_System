../ips/enc_buff/synth/enc_buff.vhd