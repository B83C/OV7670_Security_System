../ips/rgb_stack/synth/rgb_stack.vhd