ips/buffer_mem/synth/buffer_mem.vhd